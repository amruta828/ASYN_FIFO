`define DSIZE 8
`define no_of_transactions 16
